/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): M. Ceska, J. Matyas, V. Mrazek, and T. Vojnar,  Designing Approximate Arithmetic Circuits with Combined Error Constraints. In: Proceeding of 25th Euromicro Conference on Digital System Design 2022 (DSD'22). Gran Canaria, 2022. 
* This file contains a circuit from a sub-set of pareto optimal circuits with respect to the pwr and mre parameters
***/
// MAE% = 0.44 %
// MAE = 285 
// WCE% = 4.13 %
// WCE = 2709 
// WCRE% = 125.00 %
// EP% = 98.68 %
// MRE% = 5.03 %
// MSE = 172520 
// PDK45_PWR = 0.142 mW
// PDK45_AREA = 347.8 um2
// PDK45_DELAY = 0.91 ns

module mul8u_2NDH (
	A,
	B,
	Z
);

input [7:0] A;
input [7:0] B;
output [15:0] O;

wire sig_18;
wire sig_20;
wire sig_21;
wire sig_23;
wire sig_24;
wire sig_27;
wire sig_31;
wire sig_33;
wire sig_36;
wire sig_37;
wire sig_39;
wire sig_42;
wire sig_43;
wire sig_44;
wire sig_45;
wire sig_49;
wire sig_50;
wire sig_51;
wire sig_52;
wire sig_53;
wire sig_54;
wire sig_55;
wire sig_56;
wire sig_58;
wire sig_59;
wire sig_60;
wire sig_63;
wire sig_64;
wire sig_65;
wire sig_69;
wire sig_73;
wire sig_78;
wire sig_79;
wire sig_81;
wire sig_84;
wire sig_86;
wire sig_91;
wire sig_92;
wire sig_93;
wire sig_94;
wire sig_99;
wire sig_100;
wire sig_103;
wire sig_104;
wire sig_112;
wire sig_116;
wire sig_121;
wire sig_124;
wire sig_125;
wire sig_129;
wire sig_131;
wire sig_133;
wire sig_134;
wire sig_138;
wire sig_143;
wire sig_146;
wire sig_147;
wire sig_148;
wire sig_149;
wire sig_151;
wire sig_153;
wire sig_157;
wire sig_161;
wire sig_163;
wire sig_164;
wire sig_165;
wire sig_166;
wire sig_167;
wire sig_168;
wire sig_172;
wire sig_173;
wire sig_176;
wire sig_179;
wire sig_180;
wire sig_181;
wire sig_183;
wire sig_187;
wire sig_193;
wire sig_197;
wire sig_201;
wire sig_202;
wire sig_203;
wire sig_206;
wire sig_207;
wire sig_208;
wire sig_213;
wire sig_216;
wire sig_217;
wire sig_218;
wire sig_219;
wire sig_220;
wire sig_221;
wire sig_222;
wire sig_223;
wire sig_224;
wire sig_228;
wire sig_230;
wire sig_232;
wire sig_233;
wire sig_235;
wire sig_238;
wire sig_240;
wire sig_248;
wire sig_251;
wire sig_253;
wire sig_256;
wire sig_257;
wire sig_258;
wire sig_259;
wire sig_264;
wire sig_266;
wire sig_267;
wire sig_269;
wire sig_274;
wire sig_275;
wire sig_276;
wire sig_281;
wire sig_287;
wire sig_289;
wire sig_290;
wire sig_292;
wire sig_297;
wire sig_302;
wire sig_304;
wire sig_309;
wire sig_322;
wire sig_330;
wire sig_349;
wire sig_350;
wire sig_353;
wire sig_354;
wire sig_356;
wire sig_357;
wire sig_358;
wire sig_359;
wire sig_360;
wire sig_361;
wire sig_362;

assign sig_18 = A[7] & B[5];
assign sig_20 = A[4] & B[7];
assign sig_21 = A[0] & B[7];
assign sig_23 = A[7] & B[1];
assign sig_24 = A[2] & B[5];
assign sig_27 = A[3] & B[5];
assign sig_31 = A[5] & B[7];
assign sig_33 = A[4] & B[4];
assign sig_36 = A[2] & B[6];
assign sig_37 = A[7] & B[3];
assign sig_39 = A[6] & B[4];
assign sig_42 = A[4] & B[3];
assign sig_43 = A[6] & B[2];
assign sig_44 = A[3] & B[4];
assign sig_45 = A[6] & B[6];
assign sig_49 = A[7] & B[2];
assign sig_50 = A[6] & B[3];
assign sig_51 = A[1] & B[7];
assign sig_52 = A[7] & B[0];
assign sig_53 = A[7] & B[4];
assign sig_54 = A[3] & B[6];
assign sig_55 = A[1] & B[6];
assign sig_56 = A[5] & B[6];
assign sig_58 = A[6] & B[7];
assign sig_59 = A[5] & B[2];
assign sig_60 = A[5] & B[4];
assign sig_63 = A[5] & B[5];
assign sig_64 = A[7] & B[6];
assign sig_65 = A[3] & B[7];
assign sig_69 = A[6] & B[1];
assign sig_73 = A[7] & B[7];
assign sig_78 = A[4] & B[5];
assign sig_79 = A[5] & B[3];
assign sig_81 = A[2] & B[7];
assign sig_84 = A[6] & B[5];
assign sig_86 = A[4] & B[6];
assign sig_91 = sig_23 | sig_43;
assign sig_92 = sig_58 & sig_64;
assign sig_93 = sig_64 ^ sig_58;
assign sig_94 = sig_50 | sig_60;
assign sig_99 = sig_37 ^ sig_39;
assign sig_100 = sig_37 & sig_39;
assign sig_103 = sig_99 ^ sig_63;
assign sig_104 = sig_79 | sig_33;
assign sig_112 = sig_42 | sig_36;
assign sig_116 = sig_94 | sig_78;
assign sig_121 = sig_79 & sig_39;
assign sig_124 = sig_78 & sig_94;
assign sig_125 = sig_73 ^ sig_92;
assign sig_129 = sig_84 & sig_53;
assign sig_131 = sig_53 ^ sig_84;
assign sig_133 = sig_129 ^ sig_45;
assign sig_134 = sig_31 & sig_133;
assign sig_138 = sig_63 & sig_99;
assign sig_143 = sig_24 | sig_44;
assign sig_146 = sig_100 | sig_138;
assign sig_147 = sig_143 | sig_55;
assign sig_148 = sig_104 | sig_27;
assign sig_149 = sig_124 & B[6];
assign sig_151 = sig_146 ^ sig_56;
assign sig_153 = sig_133 ^ sig_31;
assign sig_157 = sig_124 ^ sig_86;
assign sig_161 = sig_49 | sig_116;
assign sig_163 = sig_116 & sig_49;
assign sig_164 = sig_103 ^ sig_163;
assign sig_165 = sig_146 & sig_56;
assign sig_166 = sig_153 & sig_18;
assign sig_167 = sig_112 | sig_59;
assign sig_168 = sig_151 ^ sig_20;
assign sig_172 = sig_121 | sig_54;
assign sig_173 = sig_93 & sig_166;
assign sig_176 = sig_129 & B[6];
assign sig_179 = sig_131 ^ sig_168;
assign sig_180 = sig_91 ^ sig_167;
assign sig_181 = sig_168 & sig_131;
assign sig_183 = sig_157 | sig_65;
assign sig_187 = sig_103 & sig_163;
assign sig_193 = sig_20 & sig_151;
assign sig_197 = sig_18 ^ sig_153;
assign sig_201 = sig_176 | sig_134;
assign sig_202 = sig_93 ^ sig_166;
assign sig_203 = sig_65 & sig_157;
assign sig_206 = sig_165 | sig_193;
assign sig_207 = sig_91 & sig_167;
assign sig_208 = sig_197 & sig_181;
assign sig_213 = sig_164 ^ sig_183;
assign sig_216 = sig_197 ^ sig_181;
assign sig_217 = sig_201 & sig_202;
assign sig_218 = sig_149 | sig_203;
assign sig_219 = sig_148 & sig_180;
assign sig_220 = sig_36 | sig_51;
assign sig_221 = sig_173 | sig_217;
assign sig_222 = sig_202 ^ sig_201;
assign sig_223 = sig_183 & sig_164;
assign sig_224 = sig_180 ^ sig_148;
assign sig_228 = sig_73 & sig_221;
assign sig_230 = sig_206 & sig_216;
assign sig_232 = sig_216 ^ sig_206;
assign sig_233 = sig_187 | sig_223;
assign sig_235 = sig_172 | sig_81;
assign sig_238 = sig_125 ^ sig_221;
assign sig_240 = sig_179 & sig_233;
assign sig_248 = sig_208 | sig_230;
assign sig_251 = sig_207 | sig_219;
assign sig_253 = sig_179 ^ sig_233;
assign sig_256 = sig_161 ^ sig_251;
assign sig_257 = sig_222 ^ sig_248;
assign sig_258 = sig_222 & sig_248;
assign sig_259 = sig_235 & sig_256;
assign sig_264 = sig_253 ^ sig_218;
assign sig_266 = sig_218 & sig_253;
assign sig_267 = sig_240 | sig_266;
assign sig_269 = sig_161 & sig_251;
assign sig_274 = sig_256 ^ sig_235;
assign sig_275 = sig_232 & sig_267;
assign sig_276 = sig_232 ^ sig_267;
assign sig_281 = sig_222 & sig_275;
assign sig_287 = sig_269 | sig_259;
assign sig_289 = sig_224 | sig_220;
assign sig_290 = sig_147 | sig_69;
assign sig_292 = sig_258 | sig_281;
assign sig_297 = sig_290 | sig_52;
assign sig_302 = sig_213 & sig_287;
assign sig_304 = sig_213 ^ sig_287;
assign sig_309 = sig_297 | sig_21;
assign sig_322 = sig_264 ^ sig_302;
assign sig_330 = sig_264 & sig_302;
assign sig_349 = sig_276 ^ sig_330;
assign sig_350 = sig_276 & sig_330;
assign sig_353 = sig_257 & sig_350;
assign sig_354 = sig_275 | sig_350;
assign sig_356 = sig_257 ^ sig_354;
assign sig_357 = sig_292 | sig_353;
assign sig_358 = sig_238 ^ sig_357;
assign sig_359 = sig_322;
assign sig_360 = sig_73 & sig_357;
assign sig_361 = sig_228 | sig_360;
assign sig_362 = sig_92 | sig_361;

assign O[0] = sig_151;
assign O[1] = sig_222;
assign O[2] = sig_143;
assign O[3] = sig_143;
assign O[4] = sig_290;
assign O[5] = sig_289;
assign O[6] = sig_309;
assign O[7] = sig_309;
assign O[8] = sig_289;
assign O[9] = sig_274;
assign O[10] = sig_304;
assign O[11] = sig_359;
assign O[12] = sig_349;
assign O[13] = sig_356;
assign O[14] = sig_358;
assign O[15] = sig_362;

endmodule



